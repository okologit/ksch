//========================================================================================================================
// UART SELECTOR
//========================================================================================================================


module uart_selector

#(parameter CHANNEL_AMOUNT = 8)

//========================================================================================================================

(
input clk, reset, en,
input [15:0] d_bus,

output logic [CHANNEL_AMOUNT-1:0] uart_en
);

//========================================================================================================================

logic [1:0] en_sync;
logic [1:0] [15:0] d_bus_sync;

//========================================================================================================================

always_ff @ (posedge clk or posedge reset) begin

  en_sync <= {en_sync[0], en};
  d_bus_sync <= {d_bus_sync[0], d_bus};

  if (reset)
     uart_en <= 'd0;
  else if (en_sync[1])
     case (d_bus_sync[1])
           'd1, 'd2, 'd4, 'd8, 'd16, 'd32, 'd64, 'd128 :
              uart_en <= d_bus_sync[1][CHANNEL_AMOUNT-1:0];
     default: uart_en <= 'd0;
     endcase
  else
     uart_en <= 'd0;

end


endmodule
